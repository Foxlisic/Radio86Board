module vg75
(
    input           clock,
    output          r,
    output          g,
    output          b,
    output          hs,
    output          vs
);

endmodule
